magic
tech sky130A
magscale 1 2
timestamp 1734384604
<< checkpaint >>
rect -1556 -1539 1556 1539
<< pwell >>
rect -296 -279 296 279
<< nmos >>
rect -100 -131 100 69
<< ndiff >>
rect -158 57 -100 69
rect -158 -119 -146 57
rect -112 -119 -100 57
rect -158 -131 -100 -119
rect 100 57 158 69
rect 100 -119 112 57
rect 146 -119 158 57
rect 100 -131 158 -119
<< ndiffc >>
rect -146 -119 -112 57
rect 112 -119 146 57
<< psubdiff >>
rect -260 209 260 243
rect -260 -209 -226 209
rect 226 -209 260 209
rect -260 -243 -164 -209
rect 164 -243 260 -209
<< psubdiffcont >>
rect -164 -243 164 -209
<< poly >>
rect -100 141 100 157
rect -100 107 -84 141
rect 84 107 100 141
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -84 107 84 141
<< locali >>
rect -260 209 260 243
rect -260 -209 -226 209
rect -100 107 -84 141
rect 84 107 100 141
rect -146 57 -112 73
rect -146 -135 -112 -119
rect 112 57 146 73
rect 112 -135 146 -119
rect 226 -209 260 209
rect -260 -243 -164 -209
rect 164 -243 260 -209
<< properties >>
string FIXED_BBOX -243 -226 243 226
<< end >>
