magic
tech sky130A
magscale 1 2
timestamp 1734384604
<< checkpaint >>
rect -1556 -1644 1556 1644
<< nwell >>
rect -296 -384 296 384
<< pmos >>
rect -100 -236 100 164
<< pdiff >>
rect -158 152 -100 164
rect -158 -224 -146 152
rect -112 -224 -100 152
rect -158 -236 -100 -224
rect 100 152 158 164
rect 100 -224 112 152
rect 146 -224 158 152
rect 100 -236 158 -224
<< pdiffc >>
rect -146 -224 -112 152
rect 112 -224 146 152
<< nsubdiff >>
rect -260 314 260 348
rect -260 -314 -226 314
rect 226 -314 260 314
rect -260 -348 -164 -314
rect 164 -348 260 -314
<< nsubdiffcont >>
rect -164 -348 164 -314
<< poly >>
rect -100 245 100 261
rect -100 211 -84 245
rect 84 211 100 245
rect -100 164 100 211
rect -100 -262 100 -236
<< polycont >>
rect -84 211 84 245
<< locali >>
rect -260 314 260 348
rect -260 -314 -226 314
rect -100 211 -84 245
rect 84 211 100 245
rect -146 152 -112 168
rect -146 -240 -112 -224
rect 112 152 146 168
rect 112 -240 146 -224
rect 226 -314 260 314
rect -260 -348 -164 -314
rect 164 -348 260 -314
<< properties >>
string FIXED_BBOX -243 -331 243 331
<< end >>
