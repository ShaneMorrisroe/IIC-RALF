magic
tech sky130A
magscale 1 2
timestamp 1734384604
<< checkpaint >>
rect 181 2336 3259 2436
rect 181 1656 5143 2336
rect -1539 1644 5143 1656
rect -1556 1556 5143 1644
rect -1644 1539 5143 1556
rect -1656 -876 5143 1539
rect -1656 -1539 1656 -876
rect 1855 -1368 5143 -876
rect -1644 -1556 1644 -1539
rect -1556 -1644 1556 -1556
rect -1539 -1656 1539 -1644
use XM1  XM1_0 ~/IIC-RALF/Magic/Devices
timestamp 1734384604
transform 0 1 2278 -1 0 780
box -296 -279 296 279
use XM2  XM2_0 ~/IIC-RALF/Magic/Devices
timestamp 1734384604
transform 0 1 2836 -1 0 780
box -296 -279 296 279
use XM3  XM3_0 ~/IIC-RALF/Magic/Devices
timestamp 1734384604
transform 0 1 3499 -1 0 780
box -296 -384 296 384
use XM4  XM4_0 ~/IIC-RALF/Magic/Devices
timestamp 1734384604
transform 0 1 3499 -1 0 188
box -296 -384 296 384
use XM5  XM5_0 ~/IIC-RALF/Magic/Devices
timestamp 1734384604
transform 0 1 1720 -1 0 780
box -396 -279 396 279
<< end >>
